`include "top.sv"